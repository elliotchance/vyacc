module main

// FILE *fopen(const char *file_name, const char *mode_of_operation)
// fn fopen(file_name string, mode_of_operation string) ?os.File {
// 	return os.open_file(file_name, mode_of_operation) or {
// 		return none
// 	}
// }

// int fprintf(FILE *stream, const char *format, ...)
// fn fprintf(stream os.File, format string, ...) int {
// 	return 0
// }
