module main

// defines for constructing filenames

const code_suffix = '.code.v'
const defines_suffix = '.tab.h.v' // If this is removed, update README
const output_suffix = '.tab.v'
const verbose_suffix = '.output'
